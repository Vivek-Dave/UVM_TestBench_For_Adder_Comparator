
`include "interface.sv"
`include "tb_pkg.sv"
module top;
  import uvm_pkg::*;
  import tb_pkg::*;
  
  //----------------------------------------------------------------------------
  intf i_intf();
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  add_comp DUT(.n1(i_intf.n1),
               .n2(i_intf.n2),
               .enabel_sum(i_intf.enabel_sum),
               .sum(i_intf.sum),
               .more(i_intf.more),
               .less(i_intf.less),
               .match(i_intf.match)
               );
  //----------------------------------------------------------------------------               
 
  //----------------------------------------------------------------------------
  initial begin
    $dumpfile("dumpfile.vcd");
    $dumpvars;
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    uvm_config_db#(virtual intf)::set(uvm_root::get(),"","vif",i_intf);
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    run_test("add_comp_test");
  end
  //----------------------------------------------------------------------------
endmodule

