
interface intf();
    // ------------------- port declaration-------------------------------------
    logic [7:0]   n1;
    logic [7:0]   n2;
    logic enabel_sum;
    logic [8:0]  sum;
    logic       more;
    logic       less;
    logic      match;
    //--------------------------------------------------------------------------

endinterface

